interface encoder_if(input logic clk, input logic reset);
    // Define interface signals
    logic [3:0] in_data;
    logic [1:0] out_data;
endinterface
